package instructions is
	constant halt : std_logic_vector := "111111";
	constant nop : std_logic_vector := "000000";
	constant load_reg_reg : std_logic_vector := "000001";
	constant load8_reg_reg : std_logic_vector := "000010";
	constant load_reg_addr : std_logic_vector := "000011";
	constant load8_reg_addr : std_logic_vector := "000100";
	constant load-imm_reg_imm : std_logic_vector := "000101";
	constant load-addr_reg_addr : std_logic_vector := "000110";
	constant store_reg_reg : std_logic_vector := "000111";
	constant store<_reg_reg : std_logic_vector := "001000";
	constant store>_reg_reg : std_logic_vector := "001001";
	constant store_reg_addr : std_logic_vector := "001010";
	constant store<_reg_addr : std_logic_vector := "001011";
	constant store>_reg_addr : std_logic_vector := "001100";
	constant push_reg : std_logic_vector := "001101";
	constant pop_reg : std_logic_vector := "001110";
	constant add_reg_reg : std_logic_vector := "001111";
	constant sub_reg_reg : std_logic_vector := "010000";
	constant cmp_reg_reg : std_logic_vector := "010001";
	constant not_reg : std_logic_vector := "010010";
	constant shiftl_reg : std_logic_vector := "010011";
	constant shiftr_reg : std_logic_vector := "010100";
	constant and_reg_reg : std_logic_vector := "010101";
	constant or_reg_reg : std_logic_vector := "010110";
	constant xor_reg_reg : std_logic_vector := "010111";
	constant jump_addr : std_logic_vector := "011000";
	constant jump==_addr : std_logic_vector := "011001";
	constant jump<_addr : std_logic_vector := "011010";
	constant jump>_addr : std_logic_vector := "011011";
	constant jumpc_addr : std_logic_vector := "011100";
	constant in_reg_dev : std_logic_vector := "011101";
	constant out_reg_dev : std_logic_vector := "011110";
end package instructions;